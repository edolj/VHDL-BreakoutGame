----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    22:02:15 02/22/2017 
-- Design Name: 
-- Module Name:    ram32x40 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity RAM32x80 is
    Port ( clk_i 		: in  STD_LOGIC;
           addrOUT_i : in  STD_LOGIC_VECTOR (4 downto 0);
           data_o 	: out  STD_LOGIC_VECTOR (0 to 79));
end RAM32x80;

architecture Behavioral of RAM32x80 is

	type ram_type is array (29 downto 0) of std_logic_vector (0 to 79);
   signal RAM : ram_type;
	signal dataOUT : STD_LOGIC_VECTOR (0 to 79);

begin
	
	data_o <= dataOUT;

	-- to je dvokanalni RAM. Pisemo na naslov addrIN_i, istocasno lahko beremo z naslova addrOUT_i
	-- RAM ima asinhronski bralni dostop, tako da ga je easy za uporabit. Ko naslovis, takoj dobis podatke.
	-- pisalni dostop je sinhronski.
	-- Pazi LSB bit je skrajno levi, zato da se lazje 'ujema' z organizacijo zaslona!

	process(clk_i)
	begin
		if (clk_i'event and clk_i = '1') then
			-- plosca
			RAM(0)  <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(1)  <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(2)  <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(3)  <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(4)  <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(5)  <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(6)  <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(7)  <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(8)  <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(9)  <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(10) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(11) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(12) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(13) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(14) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(15) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(16) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(17) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(18) <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
			RAM(19) <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
			RAM(20) <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
			RAM(21) <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
			RAM(22) <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
			RAM(23) <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
			RAM(24) <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
			RAM(25) <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
			RAM(26) <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
			RAM(27) <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
			RAM(28) <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
		end if;
	end process;

	dataOUT <= RAM(conv_integer(addrOUT_i));


end Behavioral;

